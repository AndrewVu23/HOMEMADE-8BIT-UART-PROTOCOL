module UART(

);
endmodule